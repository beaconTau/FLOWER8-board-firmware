// serial_flash.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module serial_flash (
		input  wire       asmi_access_granted, // asmi_access_granted.asmi_access_granted
		output wire       asmi_access_request, // asmi_access_request.asmi_access_request
		input  wire [3:0] data_in,             //             data_in.data_in
		input  wire [3:0] data_oe,             //             data_oe.data_oe
		output wire [3:0] data_out,            //            data_out.data_out
		input  wire       dclk_in,             //             dclk_in.dclkin
		input  wire       ncso_in,             //             ncso_in.scein
		input  wire       noe_in               //              noe_in.noe
	);

	altera_serial_flash_loader #(
		.INTENDED_DEVICE_FAMILY  ("Cyclone V"),
		.ENHANCED_MODE           (1),
		.ENABLE_SHARED_ACCESS    ("ON"),
		.ENABLE_QUAD_SPI_SUPPORT (1),
		.NCSO_WIDTH              (1)
	) serial_flash_loader_0 (
		.dclk_in             (dclk_in),             //             dclk_in.dclkin
		.ncso_in             (ncso_in),             //             ncso_in.scein
		.data_in             (data_in),             //             data_in.data_in
		.data_oe             (data_oe),             //             data_oe.data_oe
		.noe_in              (noe_in),              //              noe_in.noe
		.asmi_access_granted (asmi_access_granted), // asmi_access_granted.asmi_access_granted
		.data_out            (data_out),            //            data_out.data_out
		.asmi_access_request (asmi_access_request)  // asmi_access_request.asmi_access_request
	);

endmodule
