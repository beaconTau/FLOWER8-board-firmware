module power_lut(clk_i, a, z);
	 input clk_i;
    input [6:0] a;
    output reg [13:0] z;

    always @(posedge clk_i) begin
        case ({a})
            7'b0000000: z <= 14'b00000000000000;
            7'b0000001: z <= 14'b00000000000001;
            7'b0000010: z <= 14'b00000000000100;
            7'b0000011: z <= 14'b00000000001001;
            7'b0000100: z <= 14'b00000000010000;
            7'b0000101: z <= 14'b00000000011001;
            7'b0000110: z <= 14'b00000000100100;
            7'b0000111: z <= 14'b00000000110001;
            7'b0001000: z <= 14'b00000001000000;
            7'b0001001: z <= 14'b00000001010001;
            7'b0001010: z <= 14'b00000001100100;
            7'b0001011: z <= 14'b00000001111001;
            7'b0001100: z <= 14'b00000010010000;
            7'b0001101: z <= 14'b00000010101001;
            7'b0001110: z <= 14'b00000011000100;
            7'b0001111: z <= 14'b00000011100001;
            7'b0010000: z <= 14'b00000100000000;
            7'b0010001: z <= 14'b00000100100001;
            7'b0010010: z <= 14'b00000101000100;
            7'b0010011: z <= 14'b00000101101001;
            7'b0010100: z <= 14'b00000110010000;
            7'b0010101: z <= 14'b00000110111001;
            7'b0010110: z <= 14'b00000111100100;
            7'b0010111: z <= 14'b00001000010001;
            7'b0011000: z <= 14'b00001001000000;
            7'b0011001: z <= 14'b00001001110001;
            7'b0011010: z <= 14'b00001010100100;
            7'b0011011: z <= 14'b00001011011001;
            7'b0011100: z <= 14'b00001100010000;
            7'b0011101: z <= 14'b00001101001001;
            7'b0011110: z <= 14'b00001110000100;
            7'b0011111: z <= 14'b00001111000001;
            7'b0100000: z <= 14'b00010000000000;
            7'b0100001: z <= 14'b00010001000001;
            7'b0100010: z <= 14'b00010010000100;
            7'b0100011: z <= 14'b00010011001001;
            7'b0100100: z <= 14'b00010100010000;
            7'b0100101: z <= 14'b00010101011001;
            7'b0100110: z <= 14'b00010110100100;
            7'b0100111: z <= 14'b00010111110001;
            7'b0101000: z <= 14'b00011001000000;
            7'b0101001: z <= 14'b00011010010001;
            7'b0101010: z <= 14'b00011011100100;
            7'b0101011: z <= 14'b00011100111001;
            7'b0101100: z <= 14'b00011110010000;
            7'b0101101: z <= 14'b00011111101001;
            7'b0101110: z <= 14'b00100001000100;
            7'b0101111: z <= 14'b00100010100001;
            7'b0110000: z <= 14'b00100100000000;
            7'b0110001: z <= 14'b00100101100001;
            7'b0110010: z <= 14'b00100111000100;
            7'b0110011: z <= 14'b00101000101001;
            7'b0110100: z <= 14'b00101010010000;
            7'b0110101: z <= 14'b00101011111001;
            7'b0110110: z <= 14'b00101101100100;
            7'b0110111: z <= 14'b00101111010001;
            7'b0111000: z <= 14'b00110001000000;
            7'b0111001: z <= 14'b00110010110001;
            7'b0111010: z <= 14'b00110100100100;
            7'b0111011: z <= 14'b00110110011001;
            7'b0111100: z <= 14'b00111000010000;
            7'b0111101: z <= 14'b00111010001001;
            7'b0111110: z <= 14'b00111100000100;
            7'b0111111: z <= 14'b00111110000001;
            7'b1000000: z <= 14'b01000000000000;
            7'b1000001: z <= 14'b00111110000001;
            7'b1000010: z <= 14'b00111100000100;
            7'b1000011: z <= 14'b00111010001001;
            7'b1000100: z <= 14'b00111000010000;
            7'b1000101: z <= 14'b00110110011001;
            7'b1000110: z <= 14'b00110100100100;
            7'b1000111: z <= 14'b00110010110001;
            7'b1001000: z <= 14'b00110001000000;
            7'b1001001: z <= 14'b00101111010001;
            7'b1001010: z <= 14'b00101101100100;
            7'b1001011: z <= 14'b00101011111001;
            7'b1001100: z <= 14'b00101010010000;
            7'b1001101: z <= 14'b00101000101001;
            7'b1001110: z <= 14'b00100111000100;
            7'b1001111: z <= 14'b00100101100001;
            7'b1010000: z <= 14'b00100100000000;
            7'b1010001: z <= 14'b00100010100001;
            7'b1010010: z <= 14'b00100001000100;
            7'b1010011: z <= 14'b00011111101001;
            7'b1010100: z <= 14'b00011110010000;
            7'b1010101: z <= 14'b00011100111001;
            7'b1010110: z <= 14'b00011011100100;
            7'b1010111: z <= 14'b00011010010001;
            7'b1011000: z <= 14'b00011001000000;
            7'b1011001: z <= 14'b00010111110001;
            7'b1011010: z <= 14'b00010110100100;
            7'b1011011: z <= 14'b00010101011001;
            7'b1011100: z <= 14'b00010100010000;
            7'b1011101: z <= 14'b00010011001001;
            7'b1011110: z <= 14'b00010010000100;
            7'b1011111: z <= 14'b00010001000001;
            7'b1100000: z <= 14'b00010000000000;
            7'b1100001: z <= 14'b00001111000001;
            7'b1100010: z <= 14'b00001110000100;
            7'b1100011: z <= 14'b00001101001001;
            7'b1100100: z <= 14'b00001100010000;
            7'b1100101: z <= 14'b00001011011001;
            7'b1100110: z <= 14'b00001010100100;
            7'b1100111: z <= 14'b00001001110001;
            7'b1101000: z <= 14'b00001001000000;
            7'b1101001: z <= 14'b00001000010001;
            7'b1101010: z <= 14'b00000111100100;
            7'b1101011: z <= 14'b00000110111001;
            7'b1101100: z <= 14'b00000110010000;
            7'b1101101: z <= 14'b00000101101001;
            7'b1101110: z <= 14'b00000101000100;
            7'b1101111: z <= 14'b00000100100001;
            7'b1110000: z <= 14'b00000100000000;
            7'b1110001: z <= 14'b00000011100001;
            7'b1110010: z <= 14'b00000011000100;
            7'b1110011: z <= 14'b00000010101001;
            7'b1110100: z <= 14'b00000010010000;
            7'b1110101: z <= 14'b00000001111001;
            7'b1110110: z <= 14'b00000001100100;
            7'b1110111: z <= 14'b00000001010001;
            7'b1111000: z <= 14'b00000001000000;
            7'b1111001: z <= 14'b00000000110001;
            7'b1111010: z <= 14'b00000000100100;
            7'b1111011: z <= 14'b00000000011001;
            7'b1111100: z <= 14'b00000000010000;
            7'b1111101: z <= 14'b00000000001001;
            7'b1111110: z <= 14'b00000000000100;
            7'b1111111: z <= 14'b00000000000001;
            default: z <= 0;
        endcase
    end
endmodule
