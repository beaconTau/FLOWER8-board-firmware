---------------------------------------------------------------------------------
-- Univ. of Chicago  
--    --KICP--
--
-- PROJECT:      RNO-G lowthresh
-- FILE:         data_manager_simple.vhd
-- AUTHOR:       e.oberla
-- EMAIL         ejo@uchicago.edu
-- DATE:         1/2021
--
-- DESCRIPTION:  control big RAMs
--
---------------------------------------------------------------------------------
--library IEEE; 
--use ieee.std_logic_1164.all;
--use ieee.std_logic_unsigned.all;
--
--use work.defs.all;
--
--entity data_manager_simple is
--Generic(
--	
--Port(
--	adc_dA_i		: in 	std_logic_vector(3 downto 0);
--	adc_dB_i		: in 	std_logic_vector(3 downto 0);
--	adc_fclk_i	: in 	std_logic; --data frame clock
--	adc_lclk_i	: in 	std_logic; --data ddr clock
--
--	rst_i			: in 	std_logic;
--	clk_i			: in 	std_logic;
--	
--	rx_fifo_rdusedw_o : out std_logic_vector(2 downto 0);
--	rx_fifo_rd_i		: in std_logic;
--	rx_adc_data_o		: out std_logic_vector(79 downto 0);
--	serdes_clk_o:	out std_logic);
--end data_manager_simple;
--
--architecture rtl of data_manager_simple is
--
--begin
--
--
--
--end rtl;