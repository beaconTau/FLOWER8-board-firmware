---------------------------------------------------------------------------------
-- Univ. of Chicago  
--    --KICP--
--
-- PROJECT:      phased-array trigger board
-- FILE:         defs.vhd
-- AUTHOR:       e.oberla
-- EMAIL         ejo@uchicago.edu
-- DATE:         1/2016
--
-- DESCRIPTION:  type defs // register mapping
--
---------------------------------------------------------------------------------

library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--////////////////////////////////////////////////////////////////
--////////////////////////////////////////////////////////////////

--////////////////////////////////////////////////////////////////
package defs is
--////////////////////////////////////////////////////////////////

--//properties for Rx data interface from ADCs:
constant define_adc_resolution			:	integer := 7; --//no. bits
constant define_word_size					:	integer := 8; --//no. bits, size of each sample in the data array
constant define_serdes_factor 			: 	integer := 8;
constant define_adc_data_width			: 	integer := 28; 
constant define_deser_data_width			: 	integer := define_serdes_factor*define_adc_data_width;
constant pdat_size							:  integer := 2*define_serdes_factor*define_word_size; --//parallel data chunk size

--//waveform acq RAM:
constant define_ram_width  				: 	integer := 128;
constant define_ram_depth					: 	integer := 3; --// words for Rx receiving RAM (was 5 before 2/19/2018)
constant define_data_ram_depth			: 	integer := 8; --// words for block RAM -- sets time window for triggered and saved event
constant define_num_wfm_buffers			:	integer := 4; --// number of independent buffers for event waveform data

--//firmware registers:
constant define_address_size				:	integer := 8; --//8 bits for now
constant define_register_size				:	integer := 32;

--//
type adc_output_data_type is array (3 downto 0) of std_logic_vector(define_adc_data_width-1 downto 0);
type full_data_type	is array	(7 downto 0) of std_logic_vector(define_ram_width-1 downto 0);	
type RAM_CHUNKED_DATA_TYPE is array(1 downto 0) of std_logic_vector(31 downto 0);
type full_address_type	is array	(7 downto 0) of std_logic_vector(define_ram_depth-1 downto 0);	
type half_address_type  is array	(3 downto 0) of std_logic_vector(define_ram_depth-1 downto 0);	
type two_chan_address_type is array	(1 downto 0) of std_logic_vector(define_ram_depth-1 downto 0);
type full_data_address_type	is array	(7 downto 0) of std_logic_vector(define_data_ram_depth-1 downto 0);	
type aux_data_link_type is array (1 downto 0) of std_logic_vector(7 downto 0);
--//
constant surface_channels : integer := 6;
type surface_data_type is array (surface_channels-1 downto 0) of std_logic_vector(define_ram_width-1 downto 0);

--//

type event_metadata_type is array(24 downto 0) of std_logic_vector(23 downto 0);

type rx_data_delay_type is array (7 downto 0) of std_logic_vector(3 downto 0); --//delay range for rx data to align ADCs
type buffered_data_type is array (7 downto 0) of std_logic_vector(2*define_ram_width-1 downto 0);

--//registers
type register_array_type is array (2**define_address_size-1 downto 0) 
	of std_logic_vector(define_register_size-define_address_size-1 downto 0); --//8 bit address, 24 bit data

--//////////////////////////////
--//stuff for beamforming
--constant define_wave2beam_bits 	: integer := 5; --// bits involved in beamforming
--constant define_wave2beam_lo_bit : integer := 0; --// low bit from sliced adc data
--constant define_wave2beam_hi_bit : integer := define_wave2beam_lo_bit + define_wave2beam_bits; --// high bit from sliced adc data
--constant define_beam_bits			: integer := define_wave2beam_bits+3; --//effective resolution increased by 3 bits (8 antennas)
--constant define_sign_bit			: integer := define_beam_bits;
constant num_beams 					:	integer :=20;
constant num_power_bits 			:	integer :=24;
constant phased_sum_bits 			:	integer :=11;
constant phased_sum_power_bits 	:	integer :=22;
constant power_sum_bits				:	integer :=24; --actually 25 but this fits into the io regs
constant input_power_thesh_bits	:	integer :=12;

constant streaming_buffer_length	:	integer :=92;
constant phased_sum_length			:	integer :=8;
constant num_channels				:	integer :=6;

constant power_length: integer:=12;
constant power_low_bit: integer:=12;
constant power_high_bit: integer:=power_low_bit+power_length-1;



type antenna_delays is array (num_beams-1 downto 0,num_channels-1 downto 0) of integer;
constant beam_delays : antenna_delays := (others=>(others=>46));
--constant beam_delays is array (num_beams-1 down to 0) of antenna_delay :=((46,24,54,58,49,72),(46,46,46,46,46,46),others<=(0,0,0,0,0,0)); --add base offset of 46


--//data split up to samples
--type beam_data_type is array (2*define_serdes_factor*define_word_size-1 downto 0) of 
--	signed(define_beam_bits-1 downto 0);
--type beam_data_type is array (2*define_serdes_factor*define_word_size-1 downto 0) of 
--	std_logic_vector(define_beam_bits-1 downto 0);		

--constant define_num_beams : integer := 15;
--type array_of_beams_type is array (define_num_beams-1 downto 0) 
--	of std_logic_vector(2*define_serdes_factor*define_word_size-1 downto 0);
	
--////////////////////////////////
--//stuff for power detection 
--constant pow_lut_size 	: integer := 2**(define_beam_bits-1);
--constant define_pow_sum_range  : integer := 16; --//allow 16 bits

--type inst_power_array_type is array(2*define_serdes_factor-1 downto 0) of std_logic_vector(define_pow_sum_range-1 downto 0);
--type full_inst_power_array_type is array(define_num_beams-1 downto 0) of inst_power_array_type;

--type pipe_full_inst_power_array_type is array(define_num_beams-1 downto 0) of 
--	std_logic_vector(4*define_serdes_factor*define_pow_sum_range-1 downto 0);

--constant define_num_power_sums : integer := 8; --//number of sums within parallel data clock
--type sum_power_type is array(define_num_beams-1 downto 0) of 
--	std_logic_vector(define_num_power_sums*(define_pow_sum_range+1)-1 downto 0);  --//define_pos_sum_range+1 (sum of adjacent samples)
	
--/////////
--constant define_16avg_pow_sum_range : integer := 20; --//20 bits (16 bits per sample, 16 samples)
--type average_power_16samp_type is array(define_num_beams-1 downto 0) of std_logic_vector(define_16avg_pow_sum_range-1 downto 0);
----------------------------------------------------------------------
end defs;

--////////////////////////////////////////////////////////////////
--////////////////////////////////////////////////////////////////



--////////////////////////////////////////////////////////////////
package register_map is
--////////////////////////////////////////////////////////////////

constant base_adrs_dsa_cntrl		:	integer := 50;

constant base_adrs_adc_cntrl		:	integer := 54;

constant base_adrs_rdout_cntrl 	:  integer := 64;

constant base_adrs_coinc_thresh	:	integer := 86;

constant base_adrs_phased_thresh : integer :=129;
	
end register_map;
	
	
