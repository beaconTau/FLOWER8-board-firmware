
module serial_flash_loader (
	noe_in);	

	input		noe_in;
endmodule
