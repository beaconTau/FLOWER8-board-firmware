-- ChipID.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ChipID is
	port (
		clkin      : in  std_logic                     := '0'; --  clkin.clk
		reset      : in  std_logic                     := '0'; --  reset.reset
		data_valid : out std_logic;                            -- output.valid
		chip_id    : out std_logic_vector(63 downto 0)         --       .data
	);
end entity ChipID;

architecture rtl of ChipID is
	component altchip_id is
		generic (
			DEVICE_FAMILY : string                        := "";
			ID_VALUE      : std_logic_vector(63 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111"
		);
		port (
			clkin      : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			data_valid : out std_logic;                            -- valid
			chip_id    : out std_logic_vector(63 downto 0)         -- data
		);
	end component altchip_id;

begin

	chipid_inst : component altchip_id
		generic map (
			DEVICE_FAMILY => "Cyclone V",
			ID_VALUE      => "1111111111111111111111111111111111111111111111111111111111111111"
		)
		port map (
			clkin      => clkin,      --  clkin.clk
			reset      => reset,      --  reset.reset
			data_valid => data_valid, -- output.valid
			chip_id    => chip_id     --       .data
		);

end architecture rtl; -- of ChipID
