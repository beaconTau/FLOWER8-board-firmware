-- serial_flash_loader.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity serial_flash_loader is
	port (
		noe_in : in std_logic := '0'  -- noe_in.noe
	);
end entity serial_flash_loader;

architecture rtl of serial_flash_loader is
	component altera_serial_flash_loader is
		generic (
			INTENDED_DEVICE_FAMILY  : string  := "";
			ENHANCED_MODE           : boolean := true;
			ENABLE_SHARED_ACCESS    : string  := "OFF";
			ENABLE_QUAD_SPI_SUPPORT : boolean := false;
			NCSO_WIDTH              : integer := 1
		);
		port (
			noe_in : in std_logic := 'X'  -- noe
		);
	end component altera_serial_flash_loader;

begin

	serial_flash_loader_0 : component altera_serial_flash_loader
		generic map (
			INTENDED_DEVICE_FAMILY  => "Cyclone V",
			ENHANCED_MODE           => true,
			ENABLE_SHARED_ACCESS    => "OFF",
			ENABLE_QUAD_SPI_SUPPORT => true,
			NCSO_WIDTH              => 1
		)
		port map (
			noe_in => noe_in  -- noe_in.noe
		);

end architecture rtl; -- of serial_flash_loader
